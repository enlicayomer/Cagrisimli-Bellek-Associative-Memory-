library verilog;
use verilog.vl_types.all;
entity mainProject_vlg_check_tst is
    port(
        cikis0          : in     vl_logic;
        cikis1          : in     vl_logic;
        OAd0            : in     vl_logic;
        OAd1            : in     vl_logic;
        var             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mainProject_vlg_check_tst;
