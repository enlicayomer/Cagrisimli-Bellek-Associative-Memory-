library verilog;
use verilog.vl_types.all;
entity mainProject_vlg_vec_tst is
end mainProject_vlg_vec_tst;
